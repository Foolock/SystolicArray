module array16x16(
input		clk,rst,
input[15:0] a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,
input[15:0] b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15,b16,
output wire[32:0] c1,
c2, 
c3, 
c4, 
c5, 
c6, 
c7, 
c8, 
c9, 
c10, 
c11, 
c12, 
c13, 
c14, 
c15, 
c16, 
c17,
c18,
c19,
c20,
c21,
c22,
c23,
c24,
c25,
c26,
c27,
c28,
c29,
c30,
c31,
c32,
c33,
c34,
c35,
c36,
c37,
c38,
c39,
c40,
c41,
c42,
c43,
c44,
c45,
c46,
c47,
c48,
c49,
c50,
c51,
c52,
c53,
c54,
c55,
c56,
c57,
c58,
c59,
c60,
c61,
c62,
c63,
c64,
c65,
c66,
c67,
c68,
c69,
c70,
c71,
c72,
c73,
c74,
c75,
c76,
c77,
c78,
c79,
c80,
c81,
c82,
c83,
c84,
c85,
c86,
c87,
c88,
c89,
c90,
c91,
c92,
c93,
c94,
c95,
c96,
c97,
c98,
c99,
c100,
c101,
c102,
c103,
c104,
c105,
c106,
c107,
c108,
c109,
c110,
c111,
c112,
c113,
c114,
c115,
c116,
c117,
c118,
c119,
c120,
c121,
c122,
c123,
c124,
c125,
c126,
c127,
c128,
c129,
c130,
c131,
c132,
c133,
c134,
c135,
c136,
c137,
c138,
c139,
c140,
c141,
c142,
c143,
c144,
c145,
c146,
c147,
c148,
c149,
c150,
c151,
c152,
c153,
c154,
c155,
c156,
c157,
c158,
c159,
c160,
c161,
c162,
c163,
c164,
c165,
c166,
c167,
c168,
c169,
c170,
c171,
c172,
c173,
c174,
c175,
c176,
c177,
c178,
c179,
c180,
c181,
c182,
c183,
c184,
c185,
c186,
c187,
c188,
c189,
c190,
c191,
c192,
c193,
c194,
c195,
c196,
c197,
c198,
c199,
c200,
c201,
c202,
c203,
c204,
c205,
c206,
c207,
c208,
c209,
c210,
c211,
c212,
c213,
c214,
c215,
c216,
c217,
c218,
c219,
c220,
c221,
c222,
c223,
c224,
c225,
c226,
c227,
c228,
c229,
c230,
c231,
c232,
c233,
c234,
c235,
c236,
c237,
c238,
c239,
c240,
c241,
c242,
c243,
c244,
c245,
c246,
c247,
c248,
c249,
c250,
c251,
c252,
c253,
c254,
c255,
c256
);

//i stands data in x coordinate axis
wire[15:0]	i12a,i12b,i12c,i12d,i13a,i13b,i13c,i13d,i14a,i14b,i14c,i14d;
wire[15:0]	i22a,i22b,i22c,i22d,i23a,i23b,i23c,i23d,i24a,i24b,i24c,i24d;
wire[15:0]	i32a,i32b,i32c,i32d,i33a,i33b,i33c,i33d,i34a,i34b,i34c,i34d;
wire[15:0]	i42a,i42b,i42c,i42d,i43a,i43b,i43c,i43d,i44a,i44b,i44c,i44d;
//j stands data in y coordinate axis
wire[15:0]	j21a,j21b,j21c,j21d,j22a,j22b,j22c,j22d,j23a,j23b,j23c,j23d,j24a,j24b,j24c,j24d;
wire[15:0]	j31a,j31b,j31c,j31d,j32a,j32b,j32c,j32d,j33a,j33b,j33c,j33d,j34a,j34b,j34c,j34d;
wire[15:0]	j41a,j41b,j41c,j41d,j42a,j42b,j42c,j42d,j43a,j43b,j43c,j43d,j44a,j44b,j44c,j44d;

array4x4	u1(.clk(clk),.rst(rst),
.a1(a1),.a2(a2),.a3(a3),.a4(a4),
.b1(b1),.b2(b2),.b3(b3),.b4(b4),
.outa1(i12a),.outa2(i12b),.outa3(i12c),.outa4(i12d),
.outb1(j21a),.outb2(j21b),.outb3(j21c),.outb4(j21d),
.c1(c1),.c2(c2),.c3(c3),.c4(c4),.c5(c17),.c6(c18),.c7(c19),.c8(c20),.c9(c33),.c10(c34),.c11(c35),.c12(c36),.c13(c49),.c14(c50),.c15(c51),.c16(c52));

array4x4	u2(.clk(clk),.rst(rst),
.a1(i12a),.a2(i12b),.a3(i12c),.a4(i12d),
.b1(b5),.b2(b6),.b3(b7),.b4(b8),
.outa1(i13a),.outa2(i13b),.outa3(i13c),.outa4(i13d),
.outb1(j22a),.outb2(j22b),.outb3(j22c),.outb4(j22d),
.c1(c5),.c2(c6),.c3(c7),.c4(c8),.c5(c21),.c6(c22),.c7(c23),.c8(c24),.c9(c37),.c10(c38),.c11(c39),.c12(c40),.c13(c53),.c14(c54),.c15(c55),.c16(c56));

array4x4	u3(.clk(clk),.rst(rst),
.a1(i13a),.a2(i13b),.a3(i13c),.a4(i13d),
.b1(b9),.b2(b10),.b3(b11),.b4(b12),
.outa1(i14a),.outa2(i14b),.outa3(i14c),.outa4(i14d),
.outb1(j23a),.outb2(j23b),.outb3(j23c),.outb4(j23d),
.c1(c9),.c2(c10),.c3(c11),.c4(c12),.c5(c25),.c6(c26),.c7(c27),.c8(c28),.c9(c41),.c10(c42),.c11(c43),.c12(c44),.c13(c57),.c14(c58),.c15(c59),.c16(c60));

array4x4	u4(.clk(clk),.rst(rst),
.a1(i14a),.a2(i14b),.a3(i14c),.a4(i14d),
.b1(b13),.b2(b14),.b3(b15),.b4(b16),
.outa1(),.outa2(),.outa3(),.outa4(),
.outb1(j24a),.outb2(j24b),.outb3(j24c),.outb4(j24d),
.c1(c13),.c2(c14),.c3(c15),.c4(c16),.c5(c29),.c6(c30),.c7(c31),.c8(c32),.c9(c45),.c10(c46),.c11(c47),.c12(c48),.c13(c61),.c14(c62),.c15(c63),.c16(c64));

array4x4	u5(.clk(clk),.rst(rst),
.a1(a5),.a2(a6),.a3(a7),.a4(a8),
.b1(j21a),.b2(j21b),.b3(j21c),.b4(j21d),
.outa1(i22a),.outa2(i22b),.outa3(i22c),.outa4(i22d),
.outb1(j31a),.outb2(j31b),.outb3(j31c),.outb4(j31d),
.c1(c65),.c2(c66),.c3(c67),.c4(c68),.c5(c81),.c6(c82),.c7(c83),.c8(c84),.c9(c97),.c10(c98),.c11(c99),.c12(c100),.c13(c113),.c14(c114),.c15(c115),.c16(c116));

array4x4	u6(.clk(clk),.rst(rst),
.a1(i22a),.a2(i22b),.a3(i22c),.a4(i22d),
.b1(j22a),.b2(j22b),.b3(j22c),.b4(j22d),
.outa1(i23a),.outa2(i23b),.outa3(i23c),.outa4(i23d),
.outb1(j32a),.outb2(j32b),.outb3(j32c),.outb4(j32d),
.c1(c69),.c2(c70),.c3(c71),.c4(c72),.c5(c85),.c6(c86),.c7(c87),.c8(c88),.c9(c101),.c10(c102),.c11(c103),.c12(c104),.c13(c117),.c14(c118),.c15(c119),.c16(c120));

array4x4	u7(.clk(clk),.rst(rst),
.a1(i23a),.a2(i23b),.a3(i23c),.a4(i23d),
.b1(j23a),.b2(j23b),.b3(j23c),.b4(j23d),
.outa1(i24a),.outa2(i24b),.outa3(i24c),.outa4(i24d),
.outb1(j33a),.outb2(j33b),.outb3(j33c),.outb4(j33d),
.c1(c73),.c2(c74),.c3(c75),.c4(c76),.c5(c89),.c6(c90),.c7(c91),.c8(c92),.c9(c105),.c10(c106),.c11(c107),.c12(c108),.c13(c121),.c14(c122),.c15(c123),.c16(c124));

array4x4	u8(.clk(clk),.rst(rst),
.a1(i24a),.a2(i24b),.a3(i24c),.a4(i24d),
.b1(j24a),.b2(j24b),.b3(j24c),.b4(j24d),
.outa1(),.outa2(),.outa3(),.outa4(),
.outb1(j34a),.outb2(j34b),.outb3(j34c),.outb4(j34d),
.c1(c77),.c2(c78),.c3(c79),.c4(c80),.c5(c93),.c6(c94),.c7(c95),.c8(c96),.c9(c109),.c10(c110),.c11(c111),.c12(c112),.c13(c125),.c14(c126),.c15(c127),.c16(c128));

array4x4	u9(.clk(clk),.rst(rst),
.a1(a9),.a2(a10),.a3(a11),.a4(a12),
.b1(j31a),.b2(j31b),.b3(j31c),.b4(j31d),
.outa1(i32a),.outa2(i32b),.outa3(i32c),.outa4(i32d),
.outb1(j41a),.outb2(j41b),.outb3(j41c),.outb4(j41d),
.c1(c129),.c2(c130),.c3(c131),.c4(c132),.c5(c145),.c6(c146),.c7(c147),.c8(c148),.c9(c161),.c10(c162),.c11(c163),.c12(c164),.c13(c177),.c14(c178),.c15(c179),.c16(c180));

array4x4	u10(.clk(clk),.rst(rst),
.a1(i32a),.a2(i32b),.a3(i32c),.a4(i32d),
.b1(j32a),.b2(j32b),.b3(j32c),.b4(j32d),
.outa1(i33a),.outa2(i33b),.outa3(i33c),.outa4(i33d),
.outb1(j42a),.outb2(j42b),.outb3(j42c),.outb4(j42d),
.c1(c133),.c2(c134),.c3(c135),.c4(c136),.c5(c149),.c6(c150),.c7(c151),.c8(c152),.c9(c165),.c10(c166),.c11(c167),.c12(c168),.c13(c181),.c14(c182),.c15(c183),.c16(c184));

array4x4	u11(.clk(clk),.rst(rst),
.a1(i33a),.a2(i33b),.a3(i33c),.a4(i33d),
.b1(j33a),.b2(j33b),.b3(j33c),.b4(j33d),
.outa1(i34a),.outa2(i34b),.outa3(i34c),.outa4(i34d),
.outb1(j43a),.outb2(j43b),.outb3(j43c),.outb4(j43d),
.c1(c137),.c2(c138),.c3(c139),.c4(c140),.c5(c153),.c6(c154),.c7(c155),.c8(c156),.c9(c169),.c10(c170),.c11(c171),.c12(c172),.c13(c185),.c14(c186),.c15(c187),.c16(c188));

array4x4	u12(.clk(clk),.rst(rst),
.a1(i34a),.a2(i34b),.a3(i34c),.a4(i34d),
.b1(j34a),.b2(j34b),.b3(j34c),.b4(j34d),
.outa1(),.outa2(),.outa3(),.outa4(),
.outb1(j44a),.outb2(j44b),.outb3(j44c),.outb4(j44d),
.c1(c141),.c2(c142),.c3(c143),.c4(c144),.c5(c157),.c6(c158),.c7(c159),.c8(c160),.c9(c173),.c10(c174),.c11(c175),.c12(c176),.c13(c189),.c14(c190),.c15(c191),.c16(c192));

array4x4	u13(.clk(clk),.rst(rst),
.a1(a13),.a2(a14),.a3(a15),.a4(a16),
.b1(j41a),.b2(j41b),.b3(j41c),.b4(j41d),
.outa1(i42a),.outa2(i42b),.outa3(i42c),.outa4(i42d),
.outb1(),.outb2(),.outb3(),.outb4(),
.c1(c193),.c2(c194),.c3(c195),.c4(c196),.c5(c209),.c6(c210),.c7(c211),.c8(c212),.c9(c225),.c10(c226),.c11(c227),.c12(c228),.c13(c241),.c14(c242),.c15(c243),.c16(c244));

array4x4	u14(.clk(clk),.rst(rst),
.a1(i42a),.a2(i42b),.a3(i42c),.a4(i42d),
.b1(j42a),.b2(j42b),.b3(j42c),.b4(j42d),
.outa1(i43a),.outa2(i43b),.outa3(i43c),.outa4(i43d),
.outb1(),.outb2(),.outb3(),.outb4(),
.c1(c197),.c2(c198),.c3(c199),.c4(c200),.c5(c213),.c6(c214),.c7(c215),.c8(c216),.c9(c229),.c10(c230),.c11(c231),.c12(c232),.c13(c245),.c14(c246),.c15(c247),.c16(c248));

array4x4	u15(.clk(clk),.rst(rst),
.a1(i43a),.a2(i43b),.a3(i43c),.a4(i43d),
.b1(j43a),.b2(j43b),.b3(j43c),.b4(j43d),
.outa1(i44a),.outa2(i44b),.outa3(i44c),.outa4(i44d),
.outb1(),.outb2(),.outb3(),.outb4(),
.c1(c201),.c2(c202),.c3(c203),.c4(c204),.c5(c217),.c6(c218),.c7(c219),.c8(c220),.c9(c233),.c10(c234),.c11(c235),.c12(c236),.c13(c249),.c14(c250),.c15(c251),.c16(c252));

array4x4	u16(.clk(clk),.rst(rst),
.a1(i44a),.a2(i44b),.a3(i44c),.a4(i44d),
.b1(j44a),.b2(j44b),.b3(j44c),.b4(j44d),
.outa1(),.outa2(),.outa3(),.outa4(),
.outb1(),.outb2(),.outb3(),.outb4(),
.c1(c205),.c2(c206),.c3(c207),.c4(c208),.c5(c221),.c6(c222),.c7(c223),.c8(c224),.c9(c237),.c10(c238),.c11(c239),.c12(c240),.c13(c253),.c14(c254),.c15(c255),.c16(c256));

endmodule