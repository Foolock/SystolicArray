`timescale 1ns/100ps
module tb2;

reg		clk,rst;
reg[15:0] a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16;
reg[15:0] b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15,b16;
wire[32:0] c1,
c2, 
c3, 
c4, 
c5, 
c6, 
c7, 
c8, 
c9, 
c10, 
c11, 
c12, 
c13, 
c14, 
c15, 
c16, 
c17,
c18,
c19,
c20,
c21,
c22,
c23,
c24,
c25,
c26,
c27,
c28,
c29,
c30,
c31,
c32,
c33,
c34,
c35,
c36,
c37,
c38,
c39,
c40,
c41,
c42,
c43,
c44,
c45,
c46,
c47,
c48,
c49,
c50,
c51,
c52,
c53,
c54,
c55,
c56,
c57,
c58,
c59,
c60,
c61,
c62,
c63,
c64,
c65,
c66,
c67,
c68,
c69,
c70,
c71,
c72,
c73,
c74,
c75,
c76,
c77,
c78,
c79,
c80,
c81,
c82,
c83,
c84,
c85,
c86,
c87,
c88,
c89,
c90,
c91,
c92,
c93,
c94,
c95,
c96,
c97,
c98,
c99,
c100,
c101,
c102,
c103,
c104,
c105,
c106,
c107,
c108,
c109,
c110,
c111,
c112,
c113,
c114,
c115,
c116,
c117,
c118,
c119,
c120,
c121,
c122,
c123,
c124,
c125,
c126,
c127,
c128,
c129,
c130,
c131,
c132,
c133,
c134,
c135,
c136,
c137,
c138,
c139,
c140,
c141,
c142,
c143,
c144,
c145,
c146,
c147,
c148,
c149,
c150,
c151,
c152,
c153,
c154,
c155,
c156,
c157,
c158,
c159,
c160,
c161,
c162,
c163,
c164,
c165,
c166,
c167,
c168,
c169,
c170,
c171,
c172,
c173,
c174,
c175,
c176,
c177,
c178,
c179,
c180,
c181,
c182,
c183,
c184,
c185,
c186,
c187,
c188,
c189,
c190,
c191,
c192,
c193,
c194,
c195,
c196,
c197,
c198,
c199,
c200,
c201,
c202,
c203,
c204,
c205,
c206,
c207,
c208,
c209,
c210,
c211,
c212,
c213,
c214,
c215,
c216,
c217,
c218,
c219,
c220,
c221,
c222,
c223,
c224,
c225,
c226,
c227,
c228,
c229,
c230,
c231,
c232,
c233,
c234,
c235,
c236,
c237,
c238,
c239,
c240,
c241,
c242,
c243,
c244,
c245,
c246,
c247,
c248,
c249,
c250,
c251,
c252,
c253,
c254,
c255,
c256;

array16x16 uut(
.clk(clk),.rst(rst),
.a1(a1),.a2(a2),.a3(a3),.a4(a4),.a5(a5),.a6(a6),.a7(a7),.a8(a8),.a9(a9),.a10(a10),.a11(a11),.a12(a12),.a13(a13),.a14(a14),.a15(a15),.a16(a16),
.b1(b1),.b2(b2),.b3(b3),.b4(b4),.b5(b5),.b6(b6),.b7(b7),.b8(b8),.b9(b9),.b10(b10),.b11(b11),.b12(b12),.b13(b13),.b14(b14),.b15(b15),.b16(b16),
.c1(c1),
.c2(c2), 
.c3(c3), 
.c4(c4), 
.c5(c5), 
.c6(c6), 
.c7(c7), 
.c8(c8), 
.c9(c9), 
.c10(c10), 
.c11(c11), 
.c12(c12), 
.c13(c13), 
.c14(c14), 
.c15(c15), 
.c16(c16), 
.c17(c17),
.c18(c18),
.c19(c19),
.c20(c20),
.c21(c21),
.c22(c22),
.c23(c23),
.c24(c24),
.c25(c25),
.c26(c26),
.c27(c27),
.c28(c28),
.c29(c29),
.c30(c30),
.c31(c31),
.c32(c32),
.c33(c33),
.c34(c34),
.c35(c35),
.c36(c36),
.c37(c37),
.c38(c38),
.c39(c39),
.c40(c40),
.c41(c41),
.c42(c42),
.c43(c43),
.c44(c44),
.c45(c45),
.c46(c46),
.c47(c47),
.c48(c48),
.c49(c49),
.c50(c50),
.c51(c51),
.c52(c52),
.c53(c53),
.c54(c54),
.c55(c55),
.c56(c56),
.c57(c57),
.c58(c58),
.c59(c59),
.c60(c60),
.c61(c61),
.c62(c62),
.c63(c63),
.c64(c64),
.c65(c65),
.c66(c66),
.c67(c67),
.c68(c68),
.c69(c69),
.c70(c70),
.c71(c71),
.c72(c72),
.c73(c73),
.c74(c74),
.c75(c75),
.c76(c76),
.c77(c77),
.c78(c78),
.c79(c79),
.c80(c80),
.c81(c81),
.c82(c82),
.c83(c83),
.c84(c84),
.c85(c85),
.c86(c86),
.c87(c87),
.c88(c88),
.c89(c89),
.c90(c90),
.c91(c91),
.c92(c92),
.c93(c93),
.c94(c94),
.c95(c95),
.c96(c96),
.c97(c97),
.c98(c98),
.c99(c99),
.c100(c100),
.c101(c101),
.c102(c102),
.c103(c103),
.c104(c104),
.c105(c105),
.c106(c106),
.c107(c107),
.c108(c108),
.c109(c109),
.c110(c110),
.c111(c111),
.c112(c112),
.c113(c113),
.c114(c114),
.c115(c115),
.c116(c116),
.c117(c117),
.c118(c118),
.c119(c119),
.c120(c120),
.c121(c121),
.c122(c122),
.c123(c123),
.c124(c124),
.c125(c125),
.c126(c126),
.c127(c127),
.c128(c128),
.c129(c129),
.c130(c130),
.c131(c131),
.c132(c132),
.c133(c133),
.c134(c134),
.c135(c135),
.c136(c136),
.c137(c137),
.c138(c138),
.c139(c139),
.c140(c140),
.c141(c141),
.c142(c142),
.c143(c143),
.c144(c144),
.c145(c145),
.c146(c146),
.c147(c147),
.c148(c148),
.c149(c149),
.c150(c150),
.c151(c151),
.c152(c152),
.c153(c153),
.c154(c154),
.c155(c155),
.c156(c156),
.c157(c157),
.c158(c158),
.c159(c159),
.c160(c160),
.c161(c161),
.c162(c162),
.c163(c163),
.c164(c164),
.c165(c165),
.c166(c166),
.c167(c167),
.c168(c168),
.c169(c169),
.c170(c170),
.c171(c171),
.c172(c172),
.c173(c173),
.c174(c174),
.c175(c175),
.c176(c176),
.c177(c177),
.c178(c178),
.c179(c179),
.c180(c180),
.c181(c181),
.c182(c182),
.c183(c183),
.c184(c184),
.c185(c185),
.c186(c186),
.c187(c187),
.c188(c188),
.c189(c189),
.c190(c190),
.c191(c191),
.c192(c192),
.c193(c193),
.c194(c194),
.c195(c195),
.c196(c196),
.c197(c197),
.c198(c198),
.c199(c199),
.c200(c200),
.c201(c201),
.c202(c202),
.c203(c203),
.c204(c204),
.c205(c205),
.c206(c206),
.c207(c207),
.c208(c208),
.c209(c209),
.c210(c210),
.c211(c211),
.c212(c212),
.c213(c213),
.c214(c214),
.c215(c215),
.c216(c216),
.c217(c217),
.c218(c218),
.c219(c219),
.c220(c220),
.c221(c221),
.c222(c222),
.c223(c223),
.c224(c224),
.c225(c225),
.c226(c226),
.c227(c227),
.c228(c228),
.c229(c229),
.c230(c230),
.c231(c231),
.c232(c232),
.c233(c233),
.c234(c234),
.c235(c235),
.c236(c236),
.c237(c237),
.c238(c238),
.c239(c239),
.c240(c240),
.c241(c241),
.c242(c242),
.c243(c243),
.c244(c244),
.c245(c245),
.c246(c246),
.c247(c247),
.c248(c248),
.c249(c249),
.c250(c250),
.c251(c251),
.c252(c252),
.c253(c253),
.c254(c254),
.c255(c255),
.c256(c256)
);

initial begin
	rst = 0;
	#25 rst = 1;
end

initial begin
	clk = 0;
	forever #25 clk = ~clk;
end

initial begin
	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//1
	#50	a1=1; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//2
	#50	a1=2; a2=17; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//3
	#50	a1=3; a2=18; a3=1; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//4
	#50	a1=4; a2=19; a3=2; a4=17; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//5
	#50	a1=5; a2=20; a3=3; a4=18; a5=1; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//6
	#50	a1=6; a2=21; a3=4; a4=19; a5=2; a6=17; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//7
	#50	a1=7; a2=22; a3=5; a4=20; a5=3; a6=18; a7=1; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//8
	#50	a1=8; a2=23; a3=6; a4=21; a5=4; a6=19; a7=2; a8=17; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//9
	#50	a1=9; a2=24; a3=7; a4=22; a5=5; a6=20; a7=3; a8=18; a9=1; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//10
	#50	a1=10; a2=25; a3=8; a4=23; a5=6; a6=21; a7=4; a8=19; a9=2; a10=17; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;	//11
	#50	a1=11; a2=26; a3=9; a4=24; a5=7; a6=22; a7=5; a8=20; a9=3; a10=18; a11=1; a12=0; a13=0; a14=0; a15=0; a16=0;	//12
	#50	a1=12; a2=27; a3=10; a4=25; a5=8; a6=23; a7=6; a8=21; a9=4; a10=19; a11=2; a12=17; a13=0; a14=0; a15=0; a16=0;	//13
	#50	a1=13; a2=28; a3=11; a4=26; a5=9; a6=24; a7=7; a8=22; a9=5; a10=20; a11=3; a12=18; a13=1; a14=0; a15=0; a16=0;	//14
	#50	a1=14; a2=29; a3=12; a4=27; a5=10; a6=25; a7=8; a8=23; a9=6; a10=21; a11=4; a12=19; a13=2; a14=17; a15=0; a16=0;	//15
	#50	a1=15; a2=30; a3=13; a4=28; a5=11; a6=26; a7=9; a8=24; a9=7; a10=22; a11=5; a12=20; a13=3; a14=18; a15=1; a16=0;	//16
	#50	a1=16; a2=31; a3=14; a4=29; a5=12; a6=27; a7=10; a8=25; a9=8; a10=23; a11=6; a12=21; a13=4; a14=19; a15=2; a16=17;	//17
	#50	a1=0; a2=32; a3=15; a4=30; a5=13; a6=28; a7=11; a8=26; a9=9; a10=24; a11=7; a12=22; a13=5; a14=20; a15=3; a16=18;	//18
	#50	a1=1; a2=0; a3=16; a4=31; a5=14; a6=29; a7=12; a8=27; a9=10; a10=25; a11=8; a12=23; a13=6; a14=21; a15=4; a16=19;	//19
	#50	a1=0; a2=0; a3=0; a4=32; a5=15; a6=30; a7=13; a8=28; a9=11; a10=26; a11=9; a12=24; a13=7; a14=22; a15=5; a16=20;	//20
	#50	a1=0; a2=0; a3=0; a4=0; a5=16; a6=31; a7=14; a8=29; a9=12; a10=27; a11=10; a12=25; a13=8; a14=23; a15=6; a16=21;	//21
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=32; a7=15; a8=30; a9=13; a10=28; a11=11; a12=26; a13=9; a14=24; a15=7; a16=22;	//22
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=16; a8=31; a9=14; a10=29; a11=12; a12=27; a13=10; a14=25; a15=8; a16=23;	//23
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=32; a9=15; a10=30; a11=13; a12=28; a13=11; a14=26; a15=9; a16=24;	//24
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=16; a10=31; a11=14; a12=29; a13=12; a14=27; a15=10; a16=25;	//25
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=32; a11=15; a12=30; a13=13; a14=28; a15=11; a16=26;	//26
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=16; a12=31; a13=14; a14=29; a15=12; a16=27;	//27
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=32; a13=15; a14=30; a15=13; a16=28;	//28
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=16; a14=31; a15=14; a16=29;	//29
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=32; a15=15; a16=30;	//30
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=16; a16=31;	//31
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=32;	//32
	#50	a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; a8=0; a9=0; a10=0; a11=0; a12=0; a13=0; a14=0; a15=0; a16=0;
end

initial begin
	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0;
	#50	b1=1; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //1
	#50	b1=1; b2=1; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //2
	#50	b1=1; b2=1; b3=1; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //3
	#50	b1=1; b2=1; b3=1; b4=1; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //4
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //5
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //6
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //7
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //8
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //9
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; //10
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; //11
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=0; b14=0; b15=0; b16=0; //12
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=0; b15=0; b16=0; //13
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=0; b16=0; //14
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=0; //15
	#50	b1=1; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //16
	#50	b1=0; b2=1; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //17
	#50	b1=0; b2=0; b3=1; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //18
	#50	b1=0; b2=0; b3=0; b4=1; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //19
	#50	b1=0; b2=0; b3=0; b4=0; b5=1; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //20
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=1; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //21
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=1; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //22
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=1; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //23
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=1; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //24
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=1; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //25
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=1; b12=1; b13=1; b14=1; b15=1; b16=1; //26
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=1; b13=1; b14=1; b15=1; b16=1; //27
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=1; b14=1; b15=1; b16=1; //28
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=1; b15=1; b16=1; //29
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=1; b16=1; //30
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=1; b16=1; //31
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=1; //32
	#50	b1=0; b2=0; b3=0; b4=0; b5=0; b6=0; b7=0; b8=0; b9=0; b10=0; b11=0; b12=0; b13=0; b14=0; b15=0; b16=0; 
end

endmodule